 module instruction_memory(
    input wire [31:0] addr,
    output reg [31:0] instr, 
    input reg clk
);

    parameter MEM_DEPTH = 30;
    reg [31:0] memory_array [0:MEM_DEPTH-1];

    initial begin
        memory_array[0] = 32'b00000000000100000000000010001011;
        memory_array[1] = 32'b00000000000100000000000010001011; 
        memory_array[2] = 32'b00000000000100000000000010001011; 
        memory_array[3] = 32'b00000000000100000000000010001101; 
        memory_array[4] = 32'b00000000000100000000000010001101; 
        memory_array[5] = 32'b00000000000100000000000010001101; 
        memory_array[6] = 32'b00000000000100000000000010001101; 
        memory_array[7] = 32'b00000000000100000000000010001101; 
        memory_array[8] = 32'b00000000000100000000000010001101; 
        memory_array[9] = 32'b00000000000100000000000010001101; 
        memory_array[10]= 32'b00000000000100000000000010001101; 
        memory_array[11] =32'b00000000000100000000000010001101; 
        memory_array[12] =32'b00000000000100000000000010001101; 
        memory_array[13] =32'b00000000000100000000000010001101; 
        memory_array[14] =32'b00000000000100000000000010001101; 
        memory_array[15] =32'b00000000000100000000000010001101; 
        memory_array[16] =32'b00000000000100000000000010001101;
        memory_array[17] =32'b00000000000100010000000110000001; 
        memory_array[18] =32'b00000000000100010000000110000001; 
        memory_array[19] =32'b00000000000100010000000110000001; 
        memory_array[20] =32'b00000000000100010000000110000001; 
        memory_array[21] =32'b00000000000100010000000110000001; 
        memory_array[22] =32'b00000000000100010000000110000001; 
        memory_array[23] =32'b00000000000100010000000110000001; 
        memory_array[24] =32'b00000000000100010000000110000001; 
        memory_array[25] =32'b00000000000100010000000110000001; 
        memory_array[26] =32'b00000000000100010000000110000001; 
        memory_array[27] =32'b00000000000100010000000110000001; 
        memory_array[28] =32'b00000000000100010000000110000001; 
        memory_array[29] =32'b00000000000100010000000110000001; 
    end

    always @(posedge clk) begin
        instr = memory_array[addr]; 
    end

endmodule