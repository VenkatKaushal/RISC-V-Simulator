module PC_Adder (
    input [31:0] pc_in,
    input enable,
    output reg [31:0] pc_out
);

    always @(posedge enable) begin
        pc_out = pc_in + 4;
    end

endmodule